`timescale 1ns / 1ps
module imm_gen
(
    input logic [31:0] pc,
    input logic [31:0]instruction,
    output logic [31:0]i_imm,
    output logic [31:0]u_imm,
    output logic [31:0]s_imm,
    output logic [31:0]sb_imm,
    output logic [31:0]uj_imm
);
always_comb
begin
	u_imm = {instruction[31:12] ,12'b0 };
	begin
	if(instruction[31]==1)
	i_imm = {20'hFFFFF, instruction[31:20]};
	else 
	i_imm = {20'd0, instruction[31:20]};
	end
	begin
	if(instruction[31]==1)
	s_imm = {20'hFFFFF,instruction[31:25],instruction[11:7]};
	else 
	s_imm = {20'd0,instruction[31:25],instruction[11:7]};
	end
	begin
	if(instruction[31]==1)
	sb_imm = {19'h7FFFF,instruction[31],instruction[7],instruction[30:25],instruction[11:8],1'b0} + pc;
	else 
	sb_imm = {19'd0,instruction[31],instruction[7],instruction[30:25],instruction[11:8],1'b0} + pc;
	end
	begin
	if(instruction[31]==1)
	uj_imm = {11'h7FF ,instruction[31],instruction[19:12],instruction[20],instruction[30:21],1'b0} + pc;
	else 
	uj_imm = {11'd0,instruction[31],instruction[19:12],instruction[20],instruction[30:21],1'b0} + pc;
	end
end
endmodule