module RF(regwrite_i,clk_i,reset_i,rs1_i,rs2_i,rd_i,wd_i,operandA_o,operandB_o,registers)
input logic regwrite_i,clk_i,reset_i,
input logic [4:0]rs1_i,
input logic [4:0]rs2_i,
input logic [4:0]rd_i,
input logic[31:0]wd_i,
output logic[31:0]operandA_o,
output logic[31:0]operandB_o,
reg [31:0] registers [0:31];

begin 
assign operandA_o = registers[rs1_i];
assign operandAB_o = registers[rs2_i];

initial begin
register[5'b0]=32'b0;
end
begin 
always @(posedge clk_i)
if (reset_i == 0)
	begin
	if( rd_i !== 0)
	begin
		if (regwrite_i !== 0) begin
		registers[rd_i] <= wd_i;
		end
		else begin
		registers[rd_i] <= wd_i;
		end

	end
	else begin
	registers[rd_i] <= 32'b0;	
	end
	end
else begin
registers[rd_i] <= 32'b0;	
end
end
endmodule: RF